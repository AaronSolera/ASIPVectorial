module FETCH_STAGE (CLK, PC_SRC, MEM_TO_REG, ALU_RESULT, READ_DATA, WD3, INSTRUCTION);

	input         CLK, PC_SRC, MEM_TO_REG;
	input  [31:0] ALU_RESULT, READ_DATA;
	output [31:0] WD3, INSTRUCTION;
	
	logic  [31:0] W_INSTRUCTION, W_RESULT, W_PC_MUX, W_PC, W_PC_PLUS;

	N_BITS_REGISTER 
		PC_REG   (CLK, CLK, 1'b0, W_PC_MUX, W_PC),
		PIPELINE (CLK, CLK, 1'b0, W_INSTRUCTION, INSTRUCTION);
		
	INSTRUCTION_MEMORY #("C:/Users/Lenovo/Desktop/ASIVP/ASIVP/code.bin")
		INS_MEM (CLK, W_PC, W_INSTRUCTION);
		
	TWO_INPUTS_N_BITS_MUX #(32) 
		MEM_MUX (ALU_RESULT, READ_DATA, MEM_TO_REG, W_RESULT),
		PC_MUX  (W_PC_PLUS, W_RESULT, PC_SRC, W_PC_MUX);
		
	N_BITS_ADDER 
		PC_ADDER (W_PC, 32'd1, W_PC_PLUS);
		
	assign WD3 = W_RESULT;

endmodule 