module ASIVP #(parameter bits = 32)();
	
endmodule
