module EXECUTE ();

endmodule 