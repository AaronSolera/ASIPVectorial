module DECODE ();


endmodule 