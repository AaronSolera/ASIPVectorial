module ASIVP ();
	
endmodule
