module DECODE_STAGE (CLK, INSTRUCTION, REG_UPDATE, REG_S_WRITE, REG_V_WRITE, WD3, WA3, R_UPDATE, PIPELINE_D);

	input          CLK, REG_UPDATE, REG_S_WRITE, REG_V_WRITE;
	input  [31:0]  INSTRUCTION;
	input  [3:0]   WD3, WA3, R_UPDATE;
	output [188:0] PIPELINE_D;
	
	logic  [16:0]  W_CONTROL;
	logic  [31:0]  W_SD1, W_SD2, W_VD1, W_VD2, W_EXTN;
	logic  [3:0]   W_SA3_MUX;
	
	N_BITS_REGISTER #(189) 
		PIPELINE (CLK, CLK, 1'b0, 
					{INSTRUCTION[29:28],W_CONTROL,INSTRUCTION[22:19],INSTRUCTION[18:15],W_SD1,W_SD2,INSTRUCTION[10:9],W_EXTN,W_VD2,W_VD1}, 
					PIPELINE_D);
		
	TWO_INPUTS_N_BITS_MUX #(4) 
		SA3_MUX (WA3, R_UPDATE, REG_UPDATE, W_SA3_MUX);
		
	N_BITS_REGISTER_BANK
		SCALAR_REG_BANK (CLK, REG_S_WRITE, INSTRUCTION[18:15], INSTRUCTION[14:11], W_SA3_MUX, WD3, W_SD1, W_SD2),
		VECTOR_REG_BANK (CLK, REG_V_WRITE, INSTRUCTION[14:11], INSTRUCTION[18:15], WA3,       WD3, W_VD2, W_VD1);
		
	EXTEND 
		EXTN (INSTRUCTION[8:0], W_EXTN);
		
	CONTROL_UNIT 
		CNTRL_UNIT (INSTRUCTION[29:23], INSTRUCTION[31:30], 
						W_CONTROL[0],  W_CONTROL[1], W_CONTROL[2],  W_CONTROL[3],  W_CONTROL[4],  W_CONTROL[6:5], W_CONTROL[7], 
						W_CONTROL[8],  W_CONTROL[9], W_CONTROL[10], W_CONTROL[11], W_CONTROL[12], W_CONTROL[13],  W_CONTROL[14], 
						W_CONTROL[15], W_CONTROL[16]);

endmodule 