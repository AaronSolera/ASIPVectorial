module ASIVP (CLK, SWITCH, IMAGE);

	input        CLK;
	input  [4:0] SWITCH;
	output [7:0] IMAGE;
	
	logic [31:0]  WD3, INSTRUCTION;
	logic [188:0] PIPELINE_D;
	logic [115:0] PIPELINE_E;
	logic [76:0]  PIPELINE_M;
	
	FETCH_STAGE 
		F (CLK, PIPELINE_M[76], PIPELINE_M[75], PIPELINE_M[63:32], PIPELINE_M[31:0], WD3, INSTRUCTION);
	DECODE_STAGE 
		D (CLK, INSTRUCTION, PIPELINE_M[72], PIPELINE_M[73], PIPELINE_M[74], WD3, PIPELINE_M[71:68], PIPELINE_M[67:64], PIPELINE_D);
	EXECUTE_STAGE 
		E (CLK, PIPELINE_D, PIPELINE_E);
	MEMORY_STAGE 
		M (CLK, PIPELINE_E, PIPELINE_M, SWITCH, IMAGE);
	
endmodule 